module RAM_TOP
(
 //�ⲿ�����ź�
 input           Clk    ,
 input           Rst    ,
 input           Ld     ,
 input           Start  ,
 input           Sliding,
 input [7:0]     Data_in,
 
 output  [6:0]    Cursor ,
 output          Empty  ,
 output          using  ,
 output          Full   ,
 
 output  [7:0]    Dout
);
//�����ź�
wire  ld_ram1               ;           
wire  start_match1          ;
wire  sliding_window_move1  ;
wire  keep_ram1             ;
wire  keep_cursor1          ;
wire  clr_ram1              ;
wire  counter1_63_1          ;
wire  counter2_63_1          ;
wire  counter3_63_1          ;
//����
parameter   DATA_width  =8 ;
parameter   DATA_num    =64;
parameter   COUNTER_max =63;
parameter   ADDR_num    =6 ;  
 
 
                             
//��������ģ��
RAM_contorl u_RAM1_contorl(
      //���������ͨ·���ź�
      .ld_ram                 (  ld_ram1               ),
	  .start_match            (  start_match1          ),
	  .sliding_window_move    (  sliding_window_move1  ),
	  .keep_ram               (  keep_ram1             ),
	  .keep_cursor            (  keep_cursor1          ),
	  .clr_ram                (  clr_ram1              ),
	  //�����ⲿ�������ź�                               
	  .Clk                    (  Clk                   ),
	  .Rst                    (  Rst                   ),
	  .LD                     (  Ld                    ),
	  .START                  (  Start                 ),
	  .SLIDING                (  Sliding               ),
	  //������������ͨ���ı�־�ź�
	  .counter1_63             (  counter1_63_1        ),
	  .counter2_63             (  counter2_63_1        ),
	  .counter3_63             (  counter3_63_1        )

);
//��������ͨ·ģ��
RAM_datapath u_RAM_datapath1 
(             
	   //�����ⲿ�������ź�
      .clk                    (   Clk                  ),          
	  .rst                    (   Rst                  ),
	  //�������Կ���ģ����ź�                       
      .ld_ram                 (   ld_ram1              ),
      .start_match            (   start_match1         ),
      .sliding_window_move    (   sliding_window_move1 ),
      .keep_ram               (   keep_ram1            ),
      .keep_cursor            (   keep_cursor1         ),
	  .clr_ram                (   clr_ram1             ),
	                                                    
	  //�����ⲿ����������                                  
	  .data_in                (   Data_in              ),
	  
      //�ֽ��������                                      
	  .dout                   (   Dout                 ),
	  
      //�����ѹ��λ���ź�                               
	  .cursor                 (   Cursor               ),
	                                                    
	  //�����������־�ź�                            
	  .counter1_63            (   counter1_63_1        ),
	  .counter2_63            (   counter2_63_1        ),
	  .counter3_63            (   counter3_63_1        ),
	                                                    
	  //�������ͨ����״̬                                  
	  .empty                  (   Empty                ),
	  .using                  (   using                ),
	  .full                   (   Full                 )		
);

endmodule